// Verilog created by ORCAD Capture

module ADC10BREAK 
 ( 
		\0 , 
		SET, 
		CONVERT );

inout	\0 , SET, CONVERT;

initial
	begin
	end

endmodule
