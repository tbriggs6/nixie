// Verilog created by ORCAD Capture

module VDC 
 ( 
		SET, 
		\0  );

inout	SET, \0 ;

initial
	begin
	end

endmodule
